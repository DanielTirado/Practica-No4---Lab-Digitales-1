module imageROM2 (
    input logic [4:0] addRom,
    output logic [31:0] dataRom
);

    // Definición de la ROM como un array de 16 entradas de 32 bits
    logic [31:0] rom [31:0];

    // Inicializar los datos directamente en el bloque initial
    initial begin
		// Diseño de un mago con túnica y bastón
		rom[0]  = 32'b00000000000000011111100000000100;
		rom[1]  = 32'b11111111000000111111110000001110;
		rom[2]  = 32'b11111111000001111111111000011111;
		rom[3]  = 32'b11111111000011100110011100001110;
		rom[4]  = 32'b11111111000011111111111100000100;
		rom[5]  = 32'b11111111000011111111111100000100;
		rom[6]  = 32'b11111111000011111111111100000100;
		rom[7]  = 32'b11111111000011111111111100000100;
		rom[8]  = 32'b11111111001111111111111110001100;
		rom[9]  = 32'b11111111111111111111111111111110;
		rom[10] = 32'b11111111111111111111111111111110;
		rom[11] = 32'b11111111111111111111111110001110;
		rom[12] = 32'b11111111000111111111111110001110;
		rom[13] = 32'b11111111000111111111111110000100;
		rom[14] = 32'b11111111000111111111111110000100;
		rom[15] = 32'b11111111000111111111111110000100;
		rom[16] = 32'b11111111000111111111111110000100;
		rom[17] = 32'b11111111000111111111111110000100;
		rom[18] = 32'b11111111000111111111111110000100;
		rom[19] = 32'b11111110000101010110101010000100;
		rom[20] = 32'b11111110000111111111111110000100;
		rom[21] = 32'b11111110000111111111111110000100;
		rom[22] = 32'b11111100000111111111111110000100;
		rom[23] = 32'b11111100000111111111111110000100;
		rom[24] = 32'b01111100000111111111111110000100;
		rom[25] = 32'b01111100000111111111111110000100;
		rom[26] = 32'b01111000000111000000001110000100;
		rom[27] = 32'b00111000000111000000001110000100;
		rom[28] = 32'b00111000000111000000001110000100;
		rom[29] = 32'b00110000000111000000001110000100;
		rom[30] = 32'b00010000001111000000001111000100;
		rom[31] = 32'b00000000111111000000001111110110;

    end

    // Asignación de la salida a partir de la dirección
    assign dataRom = rom[addRom];

endmodule