module imageROM (
    input logic [4:0] addRom,
    output logic [31:0] dataRom
);

    // Definición de la ROM como un array de 16 entradas de 32 bits
    logic [31:0] rom [31:0];

    // Inicializar los datos directamente en el bloque initial
    initial begin
		// Diseño de un mago con túnica y bastón
		rom[0]  = 32'b00100000000011111100000000000000;
		rom[1]  = 32'b01110000000111111110000011111111;
		rom[2]  = 32'b11111000001111111111000011111111;
		rom[3]  = 32'b01110000011100110011100011111111;
		rom[4]  = 32'b00100000011111111111100011111111;
		rom[5]  = 32'b00100000011111111111100011111111;
		rom[6]  = 32'b00100000011111111111100011111111;
		rom[7]  = 32'b00100000011111111111100011111111;
		rom[8]  = 32'b00110000111111111111110011111111;
		rom[9]  = 32'b01111111111111111111111111111111;
		rom[10] = 32'b01111111111111111111111111111111;
		rom[11] = 32'b01110000111111111111111111111111;
		rom[12] = 32'b01110000111111111111110011111111;
		rom[13] = 32'b00100000111111111111110011111111;
		rom[14] = 32'b00100000111111111111110011111111;
		rom[15] = 32'b00100000111111111111110011111111;
		rom[16] = 32'b00100000111111111111110011111111;
		rom[17] = 32'b00100000111111111111110011111111;
		rom[18] = 32'b00100000111111111111110011111111;
		rom[19] = 32'b00100000101010110101010001111111;
		rom[20] = 32'b00100000111111111111110001111111;
		rom[21] = 32'b00100000111111111111110001111111;
		rom[22] = 32'b00100000111111111111110001111111;
		rom[23] = 32'b00100000111111111111110000111111;
		rom[24] = 32'b00100000111111111111110000111110;
		rom[25] = 32'b00100000111111111111110000111110;
		rom[26] = 32'b00100000111000000001110000011110;
		rom[27] = 32'b00100000111000000001110000011100;
		rom[28] = 32'b00100000111000000001110000011100;
		rom[29] = 32'b00100000111000000001110000001100;
		rom[30] = 32'b00100011111000000001111000001000;
		rom[31] = 32'b01101111111000000001111110000000;
		
		


    end

    // Asignación de la salida a partir de la dirección
    assign dataRom = rom[addRom];

endmodule